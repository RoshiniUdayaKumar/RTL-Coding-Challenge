`timescale 1ns / 1ps
module logic_gates(A,B,C);
input A,B;
output C;
assign C=A^B;
endmodule
